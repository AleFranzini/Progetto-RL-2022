30 mtime=1639747843.605962435
